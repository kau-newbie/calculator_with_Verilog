module dividend(
    //곱셈 계산할 때
    
    
    
    //나눗셈 계산할 때
);



endmodule